/*------------------------------------------------------------------------------
 * File          : apb2axi_top.sv
 * Project       : APB2AXI
 * Author        : Nir Miller & Ido Oreg
 * Creation date : Nov 2, 2025
 * Description   :
 *------------------------------------------------------------------------------*/

module apb2axi_top #() ();

endmodule