/*------------------------------------------------------------------------------
 * File          : response_hanlder.sv
 * Project       : APB2AXI
 * Author        : Nir Miller & Ido Oreg
 * Creation date : Nov 2, 2025
 * Description   : Consumes Completions from the Completion FIFO, translates them into a proper APB responses.
 *------------------------------------------------------------------------------*/

module response_hanlder #() ();

endmodule